//Camila Pereira da Silva
//projeto comparador de 1 bit
//24/04/2025

module comparadorde1bit(A,B,igual, maior, menor);
	input A, B;
	output igual, maior, menor;

	assign igual = A~^B;
	assign menor = ~A & B;
	assign maior = A & ~B;



endmodule
